--
-- VHDL Architecture Kart.myTestArchitecture.rtl
--
-- Created:
--          by - axel.amand.UNKNOWN (WE7860)
--          at - 14:05:59 10.05.2022
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE rtl OF myTestArchitecture IS
BEGIN
END ARCHITECTURE rtl;

