--
-- VHDL Package Body Kart.Kart_Student
--
-- Created:
--          by - axel.amand.UNKNOWN (WE7860)
--          at - 13:03:49 23.06.2022
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
PACKAGE BODY Kart_Student IS
END Kart_Student;
