--
-- VHDL Architecture UART.serialFrameReceiver.RTL
--
-- Created:
--          by - axel.amand.UNKNOWN (WE7860)
--          at - 09:18:40 11.05.2022
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE RTL OF serialFrameReceiver IS
BEGIN
END ARCHITECTURE RTL;

